** test_ring_single_pn circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_ring_single_pn pin1 pin2
*.PININFO pin1:B pin2:B
Pring1 pin1 net1 ring_single_pn gap=0.3u radius=5.0u doping_angle=250 length_x=0.1u length_y=0.1u
Pring3 net2 net3 ring_single_pn gap=0.3u radius=5.0u doping_angle=250 length_x=0.1u length_y=0.1u
Pring5 net4 pin2 ring_single_pn gap=0.3u radius=5.0u doping_angle=250 length_x=0.1u length_y=0.1u
Pring2 net1 net2 ring_single_pn gap=0.3u radius=5.0u doping_angle=250 length_x=0.1u length_y=0.1u
Pring4 net4 net3 ring_single_pn gap=0.3u radius=5.0u doping_angle=250 length_x=0.1u length_y=0.1u
.ends
.end
