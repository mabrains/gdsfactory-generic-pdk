** test_disk_heater circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_disk_heater pin1 pin2
*.PININFO pin1:B pin2:B
Pdisk1 pin1 net1 disk_heater radius=10.0u gap=0.2u wrap_angle_deg=180.0 parity=1 heater_width=5.0u
+ heater_extent=2.0u
Pdisk2 net2 net1 disk_heater radius=10.0u gap=0.2u wrap_angle_deg=180.0 parity=1 heater_width=5.0u
+ heater_extent=2.0u
Pdisk3 net3 net2 disk_heater radius=10.0u gap=0.2u wrap_angle_deg=180.0 parity=1 heater_width=5.0u
+ heater_extent=2.0u
Pdisk4 net3 net4 disk_heater radius=10.0u gap=0.2u wrap_angle_deg=180.0 parity=1 heater_width=5.0u
+ heater_extent=2.0u
Pdisk5 pin2 net4 disk_heater radius=10.0u gap=0.2u wrap_angle_deg=180.0 parity=1 heater_width=5.0u
+ heater_extent=2.0u
.ends
.end