** general test for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_general2 pin1 pin2 pin3 pin4
*.PININFO pin1:B pin2:B pin3:B pin4:B
Pcoupler_full1 net1 net2 net4 net3 coupler_full coupling_length=40.0u dx=10.0u dy=4.8u gap=0.5u dw=0.1u
Pdbr_tapered1 net3 net5 dbr_tapered length=10.0u period=0.85 duty_cycle=0.5 w1=0.4u w2=1.0u
+ taper_length=20.0u
Pinterdigital_capacitor1 pin2 pin3 interdigital_capacitor fingers=4 finger_length=20.0u
+ finger_gap=2.0u thickness=5.0u
Pmmi1 pin1 net2 net1 mmi1x2 width=0.5u width_taper=1u length_taper=10u length_mmi=5.5u width_mmi=2.5u
+ gap_mmi=0.25u
Pring1 net4 net4 net7 ring_single_heater gap=0.2u radius=10.0u length_x=4.0u length_y=0.6u
Ppin1 net5 net6 pin3 pin2 straight_pin_slot length=500.0u via_stack_width=10.0u
+ via_stack_slab_width=10.0u via_stack_spacing=2u via_stack_slab_spacing=2.0u
Pgrating_coupler_rectangular1 net6 grating_coupler_rectangular n_periods=20 period=0.75
+ fill_factor=0.5 width_grating=11.0u length_taper=150.0u wavelength=1.55u fiber_angle=15 slab_xmin=-1.0u slab_offset=1.0u
Pmzm1 net7 pin4 mzm length_x=500u length_y=2.0u delta_length=0.0u
.ends
.end
