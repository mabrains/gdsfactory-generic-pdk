** test_grating_coupler_elliptical circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_grating_coupler_elliptical pin1 pin2
*.PININFO pin1:B pin2:B
Pgrating_coupler_elliptical1 pin1 grating_coupler_elliptical  taper_length=16.6u
+ taper_angle=40.0 wavelength=1.554u fiber_angle=15.0 grating_line_width=0.343u   n_periods=30
+ slab_xmin=-1.0u slab_offset=2.0u
Pgrating_coupler_elliptical2 pin1 grating_coupler_elliptical  taper_length=16.6u
+ taper_angle=40.0 wavelength=1.554u fiber_angle=15.0 grating_line_width=0.343u   n_periods=30
+ slab_xmin=-1.0u slab_offset=2.0u
Pgrating_coupler_elliptical3 pin1 grating_coupler_elliptical  taper_length=16.6u
+ taper_angle=40.0 wavelength=1.554u fiber_angle=15.0 grating_line_width=0.343u   n_periods=30
+ slab_xmin=-1.0u slab_offset=2.0u
Pgrating_coupler_elliptical4 pin2 grating_coupler_elliptical  taper_length=16.6u
+ taper_angle=40.0 wavelength=1.554u fiber_angle=15.0 grating_line_width=0.343u   n_periods=30
+ slab_xmin=-1.0u slab_offset=2.0u
Pgrating_coupler_elliptical5 pin2 grating_coupler_elliptical  taper_length=16.6u
+ taper_angle=40.0 wavelength=1.554u fiber_angle=15.0 grating_line_width=0.343u   n_periods=30
+ slab_xmin=-1.0u slab_offset=2.0u
Pgrating_coupler_elliptical6 pin2 grating_coupler_elliptical  taper_length=16.6u
+ taper_angle=40.0 wavelength=1.554u fiber_angle=15.0 grating_line_width=0.343u   n_periods=30
+ slab_xmin=-1.0u slab_offset=2.0u
.ends
.end
