** test_mmi2x2_with_sbend circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_mmi2x2_with_sbend pin1 pin2 pin3 pin4
*.PININFO pin1:B pin2:B pin3:B pin4:B
Pmmi1 pin1 net2 net1 pin2 mmi2x2_with_sbend
Pmmi2 net2 net4 net3 net1 mmi2x2_with_sbend
Pmmi3 net4 net5 net6 net3 mmi2x2_with_sbend
Pmmi4 net5 pin3 pin4 net6 mmi2x2_with_sbend
.ends
.end
