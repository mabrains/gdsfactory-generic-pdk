* Extracted by KLayout with GENERIC TECH LVS runset on : 21/02/2024 14:49

* cell lidar
.SUBCKT lidar
* device instance $1 r0 *1 184.66,-139.696 straight_heater_meander
P$1 \$13 \$3 \$6 \$1 straight_heater_meander heater_width=2.5e-06
* device instance $2 r0 *1 184.66,-60.696 straight_heater_meander
P$2 \$12 \$20 \$19 \$1 straight_heater_meander heater_width=2.5e-06
* device instance $3 r0 *1 184.66,10.304 straight_heater_meander
P$3 \$40 \$31 \$33 \$1 straight_heater_meander heater_width=2.5e-06
* device instance $4 r0 *1 184.66,89.304 straight_heater_meander
P$4 \$43 \$44 \$50 \$1 straight_heater_meander heater_width=2.5e-06
* device instance $5 r0 *1 89.43,-79.186 mmi1x2
P$5 \$11 \$13 \$12 mmi1x2 length_mmi=5.500000000000001e-06 width_mmi=2.5e-06
+ gap_mmi=2.5000000000000004e-07 width_taper=1.0000000000000002e-06
+ length_taper=1.0e-05
* device instance $6 r0 *1 -10.57,-4.186 mmi1x2
P$6 o_in \$11 \$27 mmi1x2 length_mmi=5.500000000000001e-06 width_mmi=2.5e-06
+ gap_mmi=2.5000000000000004e-07 width_taper=1.0000000000000002e-06
+ length_taper=1.0e-05
* device instance $7 r0 *1 89.43,70.814 mmi1x2
P$7 \$27 \$40 \$43 mmi1x2 length_mmi=5.500000000000001e-06 width_mmi=2.5e-06
+ gap_mmi=2.5000000000000004e-07 width_taper=1.0000000000000002e-06
+ length_taper=1.0e-05
* device instance $8 r0 *1 411.651,-208.961 dbr
P$8 \$3 \$2 dbr w1=4.7600000000000003e-07 w2=5.24e-07 l1=1.59e-07 l2=1.59e-07
+ n=100.0
* device instance $9 r0 *1 411.696,-56.692 dbr
P$9 \$20 \$14 dbr w1=4.7600000000000003e-07 w2=5.24e-07 l1=1.59e-07 l2=1.59e-07
+ n=100.0
* device instance $10 r0 *1 411.696,0.829 dbr
P$10 \$31 \$32 dbr w1=4.7600000000000003e-07 w2=5.24e-07 l1=1.59e-07
+ l2=1.59e-07 n=100.0
* device instance $11 r0 *1 411.651,63.518 dbr
P$11 \$44 \$41 dbr w1=4.7600000000000003e-07 w2=5.24e-07 l1=1.59e-07
+ l2=1.59e-07 n=100.0
* device instance $12 r0 *1 686.265,-150.348 grating_coupler_elliptical
P$12 \$2 \$2 grating_coupler_elliptical taper_length=1.5e-05
* device instance $13 r0 *1 595.718,-85.869 grating_coupler_elliptical
P$13 \$14 \$14 grating_coupler_elliptical taper_length=1.5e-05
* device instance $14 r0 *1 686.265,18.619 grating_coupler_elliptical
P$14 \$32 \$32 grating_coupler_elliptical taper_length=1.5e-05
* device instance $15 r0 *1 595.718,53.098 grating_coupler_elliptical
P$15 \$41 \$41 grating_coupler_elliptical taper_length=1.5e-05
.ENDS lidar
