** test_mode_converter circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_mode_converter pin1 pin2 pin3 pin4
*.PININFO pin1:B pin2:B pin3:B pin4:B
Pmode_converter1 pin2 pin1 net2 net4 mode_converter gap=0.3u length=10.0u mm_width=1.2u mc_mm_width=1.0u
+ sm_width=0.5u
Pmode_converter2 net4 net2 net3 net5 mode_converter gap=0.3u length=10.0u mm_width=1.2u mc_mm_width=1.0u
+ sm_width=0.5u
Pmode_converter3 net5 net3 net1 net6 mode_converter gap=0.3u length=10.0u mm_width=1.2u mc_mm_width=1.0u
+ sm_width=0.5u
Pmode_converter4 net6 net1 pin3 pin4 mode_converter gap=0.3u length=10.0u mm_width=1.2u mc_mm_width=1.0u
+ sm_width=0.5u
.ends
.end
