* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.SUBCKT dbr
Pdbr1 dbr1_t1 dbr1_t2 dbr w1=1u w2=1.2u l1=0.5u l2=0.6u n=10
Pdbr2 dbr2_t1 dbr2_t2 dbr w1=1.2u w2=1u l1=0.4u l2=0.6u n=5
Pdbr3 dbr3_t1 dbr3_t2 dbr w1=0.5u w2=0.7u l1=0.4u l2=0.2u n=14
.ENDS
