** test_mmi_90degree_hybrid circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_mmi_90degree_hybrid pin3 pin4 pin1 pin2
*.PININFO pin3:B pin4:B pin1:B pin2:B
Pmmi1 pin1 pin2 net4 net3 net2 net1 mmi_90degree_hybrid width=0.5u width_taper=1u length_taper=10u
+ length_mmi=5.5u width_mmi=2.5u gap_mmi=0.25u
Pmmi2 net6 net5 net1 net2 net3 net4 mmi_90degree_hybrid width=0.5u width_taper=1u length_taper=10u
+ length_mmi=5.5u width_mmi=2.5u gap_mmi=0.25u
Pmmi3 net5 net6 net7 net8 net9 net10 mmi_90degree_hybrid width=0.5u width_taper=1u length_taper=10u
+ length_mmi=5.5u width_mmi=2.5u gap_mmi=0.25u
Pmmi4 pin4 pin3 net10 net9 net8 net7 mmi_90degree_hybrid width=0.5u width_taper=1u length_taper=10u
+ length_mmi=5.5u width_mmi=2.5u gap_mmi=0.25u
.ends
.end
