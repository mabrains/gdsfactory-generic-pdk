** test_dbr circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_dbr pin2 pin1 pin3
*.PININFO pin2:B pin1:B pin3:B
Pdbr1 pin2 net1 dbr w1=0.475u l1=0.159u w2=0.525u l2=0.159u n=10
Pdbr2 net1 net2 dbr w1=0.475u l1=0.159u w2=0.525u l2=0.159u n=10
Pdbr3 pin1 net2 dbr w1=0.475u l1=0.159u w2=0.525u l2=0.159u n=10
Pdbr4 net2 net3 dbr w1=0.475u l1=0.159u w2=0.525u l2=0.159u n=10
Pdbr5 net3 pin3 dbr w1=0.475u l1=0.159u w2=0.525u l2=0.159u n=10
.ends
.end
