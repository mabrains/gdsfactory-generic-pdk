* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt coupler
Pcoupler1 c1_t1 c1_t2 c1_t3 c1_t4 coupler length=5u gap=0.25u dx=4u dy=3u
Pcoupler2 c2_t1 c2_t2 c2_t3 c2_t4 coupler length=20u gap=0.5u dx=5u dy=5u
Pcoupler3 c3_t1 c3_t2 c3_t3 c3_t4 coupler length=30u gap=1u dx=9u dy=7u
.ends
