** test_mmi1x2 circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_mmi1x2 pin1 pin3 pin2
*.PININFO pin1:B pin3:B pin2:B
Pmmi4 pin1 net1 net2 mmi1x2 width=0.5u width_taper=1u length_taper=10u length_mmi=5.5u width_mmi=2.5u
+ gap_mmi=0.25u
Pmmi1 net2 net5 net4 mmi1x2 width=0.5u width_taper=1u length_taper=10u length_mmi=5.5u width_mmi=2.5u
+ gap_mmi=0.25u
Pmmi2 net1 net6 net3 mmi1x2 width=0.5u width_taper=1u length_taper=10u length_mmi=5.5u width_mmi=2.5u
+ gap_mmi=0.25u
Pmmi5 pin2 net3 net6 mmi1x2 width=0.5u width_taper=1u length_taper=10u length_mmi=5.5u width_mmi=2.5u
+ gap_mmi=0.25u
Pmmi3 pin3 net4 net5 mmi1x2 width=0.5u width_taper=1u length_taper=10u length_mmi=5.5u width_mmi=2.5u
+ gap_mmi=0.25u
.ends
.end
