** test_coupler_adiabatic circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_coupler_adiabatic pin1 pin2 pin3 pin4
*.PININFO pin1:B pin2:B pin3:B pin4:B
Pcoupler_adiabatic1 pin1 pin2 net1 net2 coupler_adiabatic length1=20.0u length2=50.0u length3=30.0u
+ wg_sep=1.0u input_wg_sep=3.0u output_wg_sep=3.0u dw=0.1u
Pcoupler_adiabatic3 net4 net3 net6 net5 coupler_adiabatic length1=20.0u length2=50.0u length3=30.0u
+ wg_sep=1.0u input_wg_sep=3.0u output_wg_sep=3.0u dw=0.1u
Pcoupler4 net3 net4 net1 net2 coupler length=20.0u gap=0.236u dx=10u dy=4.0u
Pcdc1 pin4 pin3 net6 net5 cdc length=30.0u gap=0.5u period=0.22 duty_cycle=0.5 width_top=2.0u
+ width_bot=0.75u dx=10u dy=1.8u
.ends
.end
