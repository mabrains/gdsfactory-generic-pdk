** test_straight_pn circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_straight_pn pin1 pin2 p_pin n_pin
*.PININFO pin1:B pin2:B p_pin:B n_pin:B
Ppn1 pin1 net1 n_pin p_pin straight_pn length=1000.0u via_stack_width=10.0u via_stack_spacing=2u
Ppn2 net1 net2 n_pin p_pin straight_pn length=1000.0u via_stack_width=10.0u via_stack_spacing=2u
Ppn3 net2 net3 n_pin p_pin straight_pn length=1000.0u via_stack_width=10.0u via_stack_spacing=2u
Ppn4 net3 net4 n_pin p_pin straight_pn length=1000.0u via_stack_width=10.0u via_stack_spacing=2u
Ppn5 net4 pin2 n_pin p_pin straight_pn length=1000.0u via_stack_width=10.0u via_stack_spacing=2u
.ends
.end
