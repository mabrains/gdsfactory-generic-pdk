** test_coupler_ring circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_coupler_ring pin2 pin1 pin3 pin4
*.PININFO pin2:B pin1:B pin3:B pin4:B
Pcoupler_ring1 pin2 net1 net2 pin1 coupler_ring gap=0.2u radius=5.0u length_x=4.0u length_extension=3.0u
Pcoupler_ring3 net3 net6 net5 net4 coupler_ring gap=0.2u radius=5.0u length_x=4.0u length_extension=3.0u
Pcoupler_ring4 net6 pin4 pin3 net5 coupler_ring gap=0.2u radius=5.0u length_x=4.0u length_extension=3.0u
Pcoupler_ring2 net1 net3 net4 net2 coupler_ring gap=0.2u radius=5.0u length_x=4.0u length_extension=3.0u
.ends
.end
