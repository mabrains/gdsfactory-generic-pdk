* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt disk_simple
Pdisk1 c1_t1 c1_t2 disk raduis=8u gap=0.5u
Pdisk2 c2_t1 c2_t2 disk raduis=8u gap=0.5u
Pdisk3 c3_t1 c3_t2 disk raduis=10u gap=0.2u
Pdisk4 c4_t1 c4_t2 disk raduis=5u gap=0.4u
Pdisk5 c5_t1 c5_t2 disk raduis=10u gap=0.5u
.ends
