** test_grating_coupler_elliptical_lumerical circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_grating_coupler_elliptical_lumerical pin1 pin2
*.PININFO pin1:B pin2:B
Pgrating_coupler_elliptical_lumerical1 pin1 grating_coupler_elliptical_lumerical
+ parameters=[-2.43u, 0.1u, 0.48u] taper_angle=55.0 taper_length=12.6u fiber_angle=5.0 bias_gap=0.0u wavelength=1.554u 
+  
Pgrating_coupler_elliptical_lumerical2 pin1 grating_coupler_elliptical_lumerical
+ parameters=[-2.43u, 0.1u, 0.48u] taper_angle=55.0 taper_length=12.6u fiber_angle=5.0 bias_gap=0.0u wavelength=1.554u 
+  
Pgrating_coupler_elliptical_lumerical3 pin1 grating_coupler_elliptical_lumerical
+ parameters=[-2.43u, 0.1u, 0.48u] taper_angle=55.0 taper_length=12.6u fiber_angle=5.0 bias_gap=0.0u wavelength=1.554u 
+  
Pgrating_coupler_elliptical_lumerical4 pin2 grating_coupler_elliptical_lumerical
+ parameters=[-2.43u, 0.1u, 0.48u] taper_angle=55.0 taper_length=12.6u fiber_angle=5.0 bias_gap=0.0u wavelength=1.554u 
+  
Pgrating_coupler_elliptical_lumerical5 pin2 grating_coupler_elliptical_lumerical
+ parameters=[-2.43u, 0.1u, 0.48u] taper_angle=55.0 taper_length=12.6u fiber_angle=5.0 bias_gap=0.0u wavelength=1.554u 
+  
Pgrating_coupler_elliptical_lumerical6 pin2 grating_coupler_elliptical_lumerical
+ parameters=[-2.43u, 0.1u, 0.48u] taper_angle=55.0 taper_length=12.6u fiber_angle=5.0 bias_gap=0.0u wavelength=1.554u 
+  
.ends
.end
