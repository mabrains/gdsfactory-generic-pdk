** test_resistance_sheet circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

..subckt test_resistance_sheet pin2 pin1 pin3
*.PININFO pin2:B pin1:B pin3:B
Presistance_sheet1 pin2 net1 resistance_sheet width=10u pad_pitch=100u
Presistance_sheet2 net1 net2 resistance_sheet width=10u pad_pitch=100u
Presistance_sheet3 pin1 net2 resistance_sheet width=10u pad_pitch=100u
Presistance_sheet4 net2 net3 resistance_sheet width=10u pad_pitch=100u
Presistance_sheet5 net3 pin3 resistance_sheet width=10u pad_pitch=100u
.ends
.end

