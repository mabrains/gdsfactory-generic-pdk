** test_grating_coupler_elliptical_trenches circuit for GenericPDK
* ===================================================================================
* Copyright (c) 2024, Mabrains LLC
* Licensed under the GNU Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU Lesser General Public License
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published
* by the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: LGPL-3.0
* ===================================================================================

.subckt test_grating_coupler_elliptical_trenches pin1 pin2
*.PININFO pin1:B pin2:B
Pgrating_coupler_elliptical_trenches1 pin1 grating_coupler_elliptical_trenches  taper_length=16.6u
+ taper_angle=30.0 wavelength=1.53u fiber_angle=15.0 grating_line_width=0.343u  p_start=26
+ n_periods=30 end_straight_length=0.2u
Pgrating_coupler_elliptical_trenches2 pin1 grating_coupler_elliptical_trenches  taper_length=16.6u
+ taper_angle=30.0 wavelength=1.53u fiber_angle=15.0 grating_line_width=0.343u  p_start=26
+ n_periods=30 end_straight_length=0.2u
Pgrating_coupler_elliptical_trenches3 pin1 grating_coupler_elliptical_trenches  taper_length=16.6u
+ taper_angle=30.0 wavelength=1.53u fiber_angle=15.0 grating_line_width=0.343u  p_start=26
+ n_periods=30 end_straight_length=0.2u
Pgrating_coupler_elliptical_trenches4 pin2 grating_coupler_elliptical_trenches  taper_length=16.6u
+ taper_angle=30.0 wavelength=1.53u fiber_angle=15.0 grating_line_width=0.343u  p_start=26
+ n_periods=30 end_straight_length=0.2u
Pgrating_coupler_elliptical_trenches5 pin2 grating_coupler_elliptical_trenches  taper_length=16.6u
+ taper_angle=30.0 wavelength=1.53u fiber_angle=15.0 grating_line_width=0.343u  p_start=26
+ n_periods=30 end_straight_length=0.2u
Pgrating_coupler_elliptical_trenches6 pin2 grating_coupler_elliptical_trenches  taper_length=16.6u
+ taper_angle=30.0 wavelength=1.53u fiber_angle=15.0 grating_line_width=0.343u  p_start=26
+ n_periods=30 end_straight_length=0.2u
.ends
.end
